
module S_P (
	source,
	probe);	

	output	[63:0]	source;
	input	[63:0]	probe;
endmodule
