// unnamed.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module unnamed (
		input  wire        i_avalon_chip_select, // avalon_sdcard_slave.chipselect
		input  wire [7:0]  i_avalon_address,     //                    .address
		input  wire        i_avalon_read,        //                    .read
		input  wire        i_avalon_write,       //                    .write
		input  wire [3:0]  i_avalon_byteenable,  //                    .byteenable
		input  wire [31:0] i_avalon_writedata,   //                    .writedata
		output wire [31:0] o_avalon_readdata,    //                    .readdata
		output wire        o_avalon_waitrequest, //                    .waitrequest
		input  wire        i_clock,              //                 clk.clk
		inout  wire        b_SD_cmd,             //         conduit_end.b_SD_cmd
		inout  wire        b_SD_dat,             //                    .b_SD_dat
		inout  wire        b_SD_dat3,            //                    .b_SD_dat3
		output wire        o_SD_clock,           //                    .o_SD_clock
		input  wire        i_reset_n             //               reset.reset_n
	);

	Altera_UP_SD_Card_Avalon_Interface altera_up_sd_card_avalon_interface_0 (
		.i_avalon_chip_select (i_avalon_chip_select), // avalon_sdcard_slave.chipselect
		.i_avalon_address     (i_avalon_address),     //                    .address
		.i_avalon_read        (i_avalon_read),        //                    .read
		.i_avalon_write       (i_avalon_write),       //                    .write
		.i_avalon_byteenable  (i_avalon_byteenable),  //                    .byteenable
		.i_avalon_writedata   (i_avalon_writedata),   //                    .writedata
		.o_avalon_readdata    (o_avalon_readdata),    //                    .readdata
		.o_avalon_waitrequest (o_avalon_waitrequest), //                    .waitrequest
		.i_clock              (i_clock),              //                 clk.clk
		.i_reset_n            (i_reset_n),            //               reset.reset_n
		.b_SD_cmd             (b_SD_cmd),             //         conduit_end.export
		.b_SD_dat             (b_SD_dat),             //                    .export
		.b_SD_dat3            (b_SD_dat3),            //                    .export
		.o_SD_clock           (o_SD_clock)            //                    .export
	);

endmodule
