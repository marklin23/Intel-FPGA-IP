// i2c_master.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module i2c_master (
		input  wire        clk_clk,                    //                    clk.clk
		input  wire [3:0]  i2c_1_csr_address,          //              i2c_1_csr.address
		input  wire        i2c_1_csr_read,             //                       .read
		input  wire        i2c_1_csr_write,            //                       .write
		input  wire [31:0] i2c_1_csr_writedata,        //                       .writedata
		output wire [31:0] i2c_1_csr_readdata,         //                       .readdata
		input  wire        i2c_1_i2c_serial_sda_in,    //       i2c_1_i2c_serial.sda_in
		input  wire        i2c_1_i2c_serial_scl_in,    //                       .scl_in
		output wire        i2c_1_i2c_serial_sda_oe,    //                       .sda_oe
		output wire        i2c_1_i2c_serial_scl_oe,    //                       .scl_oe
		output wire        i2c_1_interrupt_sender_irq, // i2c_1_interrupt_sender.irq
		input  wire        reset_reset_n               //                  reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> i2c_1:rst_n

	altera_avalon_i2c #(
		.USE_AV_ST       (0),
		.FIFO_DEPTH      (32),
		.FIFO_DEPTH_LOG2 (5)
	) i2c_1 (
		.clk       (clk_clk),                         //            clock.clk
		.rst_n     (~rst_controller_reset_out_reset), //       reset_sink.reset_n
		.intr      (i2c_1_interrupt_sender_irq),      // interrupt_sender.irq
		.addr      (i2c_1_csr_address),               //              csr.address
		.read      (i2c_1_csr_read),                  //                 .read
		.write     (i2c_1_csr_write),                 //                 .write
		.writedata (i2c_1_csr_writedata),             //                 .writedata
		.readdata  (i2c_1_csr_readdata),              //                 .readdata
		.sda_in    (i2c_1_i2c_serial_sda_in),         //       i2c_serial.sda_in
		.scl_in    (i2c_1_i2c_serial_scl_in),         //                 .scl_in
		.sda_oe    (i2c_1_i2c_serial_sda_oe),         //                 .sda_oe
		.scl_oe    (i2c_1_i2c_serial_scl_oe),         //                 .scl_oe
		.src_data  (),                                //      (terminated)
		.src_valid (),                                //      (terminated)
		.src_ready (1'b0),                            //      (terminated)
		.snk_data  (16'b0000000000000000),            //      (terminated)
		.snk_valid (1'b0),                            //      (terminated)
		.snk_ready ()                                 //      (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
